1 1 0 1 0
1 2 0 1 0
1 3 0 2 0
2 8 1 3
2 9 1 3
1 6 0 1 0
1 7 0 1 0
0 10 2 1 2 1 8 
0 11 2 2 2 9 6 
2 14 1 11
2 15 1 11
0 16 2 2 2 2 14 
2 20 1 16
2 21 1 16
0 19 2 1 2 15 7 
3 22 2 0 2 10 20 
3 23 2 0 2 21 19 
